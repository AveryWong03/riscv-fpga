`default_nettype none

module pc(
    input logic clk,
    input logic [31:0] pctarget,
    input logic pcsrc,
    input logic stallf,
    output logic [31:0] pcf, pcfplus4
);

endmodule