`default_nettype none

module ex_mem_reg(
    input logic clk,
    input ex_mem d,
    output ex_mem q
);

endmodule