`default_nettype none

module alu(
    input logic [31:0] srca, srcb,
    input logic [2:0] alucontrol,
    output logic [31:0] aluresult,
    output logic zero
);

endmodule