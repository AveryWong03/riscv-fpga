`default_nettype none

module mem_wb_reg(
    input logic clk,
    input mem_wb_t d,
    output mem_wb_t q
);

endmodule