`default_nettype none

module mem_wb_reg(
    input logic clk,
    input mem_wb_t d,
    input logic [31:0] readdata_i,
    output logic [31:0] readdata_o, 
    output mem_wb_t q
);

endmodule