`default_nettype none

module if_id_reg(
    input logic clk, clr, en,
    input if_id d,
    output if_id q
);

endmodule