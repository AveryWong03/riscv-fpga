`default_nettype none

module mem_wb_reg(
    input logic clk,
    input mem_wb d,
    output mem_wb q
);

endmodule