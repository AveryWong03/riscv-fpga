`default_nettype none

module id_ex_reg(
    input logic clk, clr,
    input id_ex_t d,
    output id_ex_t q
);

endmodule