`default_nettype none

module foward_unit(
    input logic [31:0] rd1, rd2, result, aluresult, immext,
    input logic [1:0] forwarda, forwardb,
    input logic alusrc,
    output logic [31:0] srca, srcb
);

endmodule