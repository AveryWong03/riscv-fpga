`default_nettype none

module wb_stage(
    input mem_wb_t in,
    output logic regwrite,
    output logic [4:0] rd,
    output logic [31:0] result
);

endmodule