`default_nettype none

module if_stage(
    input logic clk, en,
    input logic [31:0] pcsrc, pctarget, pcplus4,
    output if_id out
);

endmodule