`default_nettype none

module id_ex_reg(
    input logic clk, clr,
    input id_ex_t d,
    input logic [31:0] rd1_i, rd2_i,
    output logic [31:0] rd1_o, rd2_o,
    output id_ex_t q
);

endmodule