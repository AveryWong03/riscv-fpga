`default_nettype none

module risc_core(  
);


endmodule