`default_nettype none

module ex_mem_reg(
    input logic clk,
    input ex_mem_t d,
    output ex_mem_t q
);

endmodule