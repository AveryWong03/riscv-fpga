`default_nettype none

module mem_stage(
    input logic clk,
    input ex_mem_t in,
    output mem_wb_t out
);

endmodule