`default_nettype none

module if_id_reg(
    input logic clk, clr, en,
    input if_id_t d,
    output if_id_t q
);

endmodule