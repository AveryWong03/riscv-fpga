`default_nettype none

module id_stage(
    input logic clk, regwrite_w,
    input if_id in,
    output id_ex out // rs1, rs2 need to be output to hazard unit
);

endmodule