`default_nettype none

module mem_stage(
    input logic clk,
    input ex_mem in,
    output mem_wb out
);

endmodule