`default_nettype none

module pc(
    input logic clk,
    input logic [31:0] pctarget,
    input logic pcsrc,
    input logic stall,
    output logic [31:0] pc, pcplus4
);

endmodule