`default_nettype none

module id_ex_reg(
    input logic clk, clr,
    input id_ex d,
    output id_ex q
);

endmodule